`timescale 1ns / 1ps

`include "axi_vip_0_exdes_generic.sv"
`include "axi_vip_0_mst_stimulus.sv"
`include "axi_vip_0_mem_basic_stimulus.sv"

module tb_slv_vip();


endmodule